module FFT32_top #(parameter WORD_SIZE = 16, parameter FRACTION = 8)
(
	input							i_clk,
	input 						i_rst,
	input       	[WORD_SIZE-1:0]     in0_re,
	input       	[WORD_SIZE-1:0]     in0_im,
	input       	[WORD_SIZE-1:0]     in1_re,
	input       	[WORD_SIZE-1:0]     in1_im,
	input       	[WORD_SIZE-1:0]     in2_re,
	input       	[WORD_SIZE-1:0]     in2_im,
	input       	[WORD_SIZE-1:0]     in3_re,
	input       	[WORD_SIZE-1:0]     in3_im,
	input       	[WORD_SIZE-1:0]     in4_re,
	input       	[WORD_SIZE-1:0]     in4_im,
	input       	[WORD_SIZE-1:0]     in5_re,
	input       	[WORD_SIZE-1:0]     in5_im,
	input       	[WORD_SIZE-1:0]     in6_re,
	input       	[WORD_SIZE-1:0]     in6_im,
	input       	[WORD_SIZE-1:0]     in7_re,
	input       	[WORD_SIZE-1:0]     in7_im,
	input       	[WORD_SIZE-1:0]     in8_re,
	input       	[WORD_SIZE-1:0]     in8_im,
	input       	[WORD_SIZE-1:0]     in9_re,
	input       	[WORD_SIZE-1:0]     in9_im,
	input       	[WORD_SIZE-1:0]     in10_re,
	input       	[WORD_SIZE-1:0]     in10_im,
	input       	[WORD_SIZE-1:0]     in11_re,
	input       	[WORD_SIZE-1:0]     in11_im,
	input       	[WORD_SIZE-1:0]     in12_re,
	input       	[WORD_SIZE-1:0]     in12_im,
	input       	[WORD_SIZE-1:0]     in13_re,
	input       	[WORD_SIZE-1:0]     in13_im,
	input       	[WORD_SIZE-1:0]     in14_re,
	input       	[WORD_SIZE-1:0]     in14_im,
	input       	[WORD_SIZE-1:0]     in15_re,
	input       	[WORD_SIZE-1:0]     in15_im,
	input       	[WORD_SIZE-1:0]     in16_re,
	input       	[WORD_SIZE-1:0]     in16_im,
	input       	[WORD_SIZE-1:0]     in17_re,
	input       	[WORD_SIZE-1:0]     in17_im,
	input       	[WORD_SIZE-1:0]     in18_re,
	input       	[WORD_SIZE-1:0]     in18_im,
	input       	[WORD_SIZE-1:0]     in19_re,
	input       	[WORD_SIZE-1:0]     in19_im,
	input       	[WORD_SIZE-1:0]     in20_re,
	input       	[WORD_SIZE-1:0]     in20_im,
	input       	[WORD_SIZE-1:0]     in21_re,
	input       	[WORD_SIZE-1:0]     in21_im,
	input       	[WORD_SIZE-1:0]     in22_re,
	input       	[WORD_SIZE-1:0]     in22_im,
	input       	[WORD_SIZE-1:0]     in23_re,
	input       	[WORD_SIZE-1:0]     in23_im,
	input       	[WORD_SIZE-1:0]     in24_re,
	input       	[WORD_SIZE-1:0]     in24_im,
	input       	[WORD_SIZE-1:0]     in25_re,
	input       	[WORD_SIZE-1:0]     in25_im,
	input       	[WORD_SIZE-1:0]     in26_re,
	input       	[WORD_SIZE-1:0]     in26_im,
	input       	[WORD_SIZE-1:0]     in27_re,
	input       	[WORD_SIZE-1:0]     in27_im,
	input       	[WORD_SIZE-1:0]     in28_re,
	input       	[WORD_SIZE-1:0]     in28_im,
	input       	[WORD_SIZE-1:0]     in29_re,
	input       	[WORD_SIZE-1:0]     in29_im,
	input       	[WORD_SIZE-1:0]     in30_re,
	input       	[WORD_SIZE-1:0]     in30_im,
	input       	[WORD_SIZE-1:0]     in31_re,
	input       	[WORD_SIZE-1:0]     in31_im,
	
	output       	[WORD_SIZE-1:0]     out0_re,
	output       	[WORD_SIZE-1:0]     out0_im,
	output       	[WORD_SIZE-1:0]     out1_re,
	output       	[WORD_SIZE-1:0]     out1_im,
	output       	[WORD_SIZE-1:0]     out2_re,
	output       	[WORD_SIZE-1:0]     out2_im,
	output       	[WORD_SIZE-1:0]     out3_re,
	output       	[WORD_SIZE-1:0]     out3_im,
	output       	[WORD_SIZE-1:0]     out4_re,
	output       	[WORD_SIZE-1:0]     out4_im,
	output       	[WORD_SIZE-1:0]     out5_re,
	output       	[WORD_SIZE-1:0]     out5_im,
	output       	[WORD_SIZE-1:0]     out6_re,
	output       	[WORD_SIZE-1:0]     out6_im,
	output       	[WORD_SIZE-1:0]     out7_re,
	output       	[WORD_SIZE-1:0]     out7_im,
	output       	[WORD_SIZE-1:0]     out8_re,
	output       	[WORD_SIZE-1:0]     out8_im,
	output       	[WORD_SIZE-1:0]     out9_re,
	output       	[WORD_SIZE-1:0]     out9_im,
	output       	[WORD_SIZE-1:0]     out10_re,
	output       	[WORD_SIZE-1:0]     out10_im,
	output       	[WORD_SIZE-1:0]     out11_re,
	output       	[WORD_SIZE-1:0]     out11_im,
	output       	[WORD_SIZE-1:0]     out12_re,
	output       	[WORD_SIZE-1:0]     out12_im,
	output       	[WORD_SIZE-1:0]     out13_re,
	output       	[WORD_SIZE-1:0]     out13_im,
	output       	[WORD_SIZE-1:0]     out14_re,
	output       	[WORD_SIZE-1:0]     out14_im,
	output       	[WORD_SIZE-1:0]     out15_re,
	output       	[WORD_SIZE-1:0]     out15_im,
	output       	[WORD_SIZE-1:0]     out16_re,
	output       	[WORD_SIZE-1:0]     out16_im,
	output       	[WORD_SIZE-1:0]     out17_re,
	output       	[WORD_SIZE-1:0]     out17_im,
	output       	[WORD_SIZE-1:0]     out18_re,
	output       	[WORD_SIZE-1:0]     out18_im,
	output       	[WORD_SIZE-1:0]     out19_re,
	output       	[WORD_SIZE-1:0]     out19_im,
	output       	[WORD_SIZE-1:0]     out20_re,
	output       	[WORD_SIZE-1:0]     out20_im,
	output       	[WORD_SIZE-1:0]     out21_re,
	output       	[WORD_SIZE-1:0]     out21_im,
	output       	[WORD_SIZE-1:0]     out22_re,
	output       	[WORD_SIZE-1:0]     out22_im,
	output       	[WORD_SIZE-1:0]     out23_re,
	output       	[WORD_SIZE-1:0]     out23_im,
	output       	[WORD_SIZE-1:0]     out24_re,
	output       	[WORD_SIZE-1:0]     out24_im,
	output       	[WORD_SIZE-1:0]     out25_re,
	output       	[WORD_SIZE-1:0]     out25_im,
	output       	[WORD_SIZE-1:0]     out26_re,
	output       	[WORD_SIZE-1:0]     out26_im,
	output       	[WORD_SIZE-1:0]     out27_re,
	output       	[WORD_SIZE-1:0]     out27_im,
	output       	[WORD_SIZE-1:0]     out28_re,
	output       	[WORD_SIZE-1:0]     out28_im,
	output       	[WORD_SIZE-1:0]     out29_re,
	output       	[WORD_SIZE-1:0]     out29_im,
	output       	[WORD_SIZE-1:0]     out30_re,
	output       	[WORD_SIZE-1:0]     out30_im,
	output       	[WORD_SIZE-1:0]     out31_re,
	output       	[WORD_SIZE-1:0]     out31_im,
	
	output 										o_FFT32_cycle_done,
	output			[1:0]						w_mux_switcher,
	output										w_address_switcher,
	output										w_FFT16_cycle_rst,
	output			[2:0]						w_STAGES,
	output										w_FFT16_cycle_done_delay
	
); 
	//wire	[1:0]					w_mux_switcher;
	//wire							w_address_switcher;
	//wire							w_FFT16_cycle_rst;
	//wire	[2:0]					w_STAGES;
	//wire 							w_FFT16_cycle_done;
	//wire 							w_FFT16_cycle_done_delay;
	
	wire	[WORD_SIZE-1:0]	FFT16_in0_re;
	wire	[WORD_SIZE-1:0]	FFT16_in0_im;
	wire	[WORD_SIZE-1:0]	FFT16_in1_re;
	wire	[WORD_SIZE-1:0]	FFT16_in1_im;
	wire	[WORD_SIZE-1:0]	FFT16_in2_re;
	wire	[WORD_SIZE-1:0]	FFT16_in2_im;
	wire	[WORD_SIZE-1:0]	FFT16_in3_re;
	wire	[WORD_SIZE-1:0]	FFT16_in3_im;
	wire	[WORD_SIZE-1:0]	FFT16_in4_re;
	wire	[WORD_SIZE-1:0]	FFT16_in4_im;
	wire	[WORD_SIZE-1:0]	FFT16_in5_re;
	wire	[WORD_SIZE-1:0]	FFT16_in5_im;
	wire	[WORD_SIZE-1:0]	FFT16_in6_re;
	wire	[WORD_SIZE-1:0]	FFT16_in6_im;
	wire	[WORD_SIZE-1:0]	FFT16_in7_re;
	wire	[WORD_SIZE-1:0]	FFT16_in7_im;
	wire	[WORD_SIZE-1:0]	FFT16_in8_re;
	wire	[WORD_SIZE-1:0]	FFT16_in8_im;
	wire	[WORD_SIZE-1:0]	FFT16_in9_re;
	wire	[WORD_SIZE-1:0]	FFT16_in9_im;
	wire	[WORD_SIZE-1:0]	FFT16_in10_re;
	wire	[WORD_SIZE-1:0]	FFT16_in10_im;
	wire	[WORD_SIZE-1:0]	FFT16_in11_re;
	wire	[WORD_SIZE-1:0]	FFT16_in11_im;
	wire	[WORD_SIZE-1:0]	FFT16_in12_re;
	wire	[WORD_SIZE-1:0]	FFT16_in12_im;
	wire	[WORD_SIZE-1:0]	FFT16_in13_re;
	wire	[WORD_SIZE-1:0]	FFT16_in13_im;
	wire	[WORD_SIZE-1:0]	FFT16_in14_re;
	wire	[WORD_SIZE-1:0]	FFT16_in14_im;
	wire	[WORD_SIZE-1:0]	FFT16_in15_re;
	wire	[WORD_SIZE-1:0]	FFT16_in15_im;
	
	wire	[WORD_SIZE-1:0]	FFT16_out0_re;
	wire	[WORD_SIZE-1:0]	FFT16_out0_im;
	wire	[WORD_SIZE-1:0]	FFT16_out1_re;
	wire	[WORD_SIZE-1:0]	FFT16_out1_im;
	wire	[WORD_SIZE-1:0]	FFT16_out2_re;
	wire	[WORD_SIZE-1:0]	FFT16_out2_im;
	wire	[WORD_SIZE-1:0]	FFT16_out3_re;
	wire	[WORD_SIZE-1:0]	FFT16_out3_im;
	wire	[WORD_SIZE-1:0]	FFT16_out4_re;
	wire	[WORD_SIZE-1:0]	FFT16_out4_im;
	wire	[WORD_SIZE-1:0]	FFT16_out5_re;
	wire	[WORD_SIZE-1:0]	FFT16_out5_im;
	wire	[WORD_SIZE-1:0]	FFT16_out6_re;
	wire	[WORD_SIZE-1:0]	FFT16_out6_im;
	wire	[WORD_SIZE-1:0]	FFT16_out7_re;
	wire	[WORD_SIZE-1:0]	FFT16_out7_im;
	wire	[WORD_SIZE-1:0]	FFT16_out8_re;
	wire	[WORD_SIZE-1:0]	FFT16_out8_im;
	wire	[WORD_SIZE-1:0]	FFT16_out9_re;
	wire	[WORD_SIZE-1:0]	FFT16_out9_im;
	wire	[WORD_SIZE-1:0]	FFT16_out10_re;
	wire	[WORD_SIZE-1:0]	FFT16_out10_im;
	wire	[WORD_SIZE-1:0]	FFT16_out11_re;
	wire	[WORD_SIZE-1:0]	FFT16_out11_im;
	wire	[WORD_SIZE-1:0]	FFT16_out12_re;
	wire	[WORD_SIZE-1:0]	FFT16_out12_im;
	wire	[WORD_SIZE-1:0]	FFT16_out13_re;
	wire	[WORD_SIZE-1:0]	FFT16_out13_im;
	wire	[WORD_SIZE-1:0]	FFT16_out14_re;
	wire	[WORD_SIZE-1:0]	FFT16_out14_im;
	wire	[WORD_SIZE-1:0]	FFT16_out15_re;
	wire	[WORD_SIZE-1:0]	FFT16_out15_im;	
	
	wire	[WORD_SIZE-1:0]	w_buffer_out0_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out0_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out1_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out1_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out2_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out2_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out3_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out3_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out4_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out4_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out5_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out5_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out6_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out6_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out7_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out7_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out8_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out8_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out9_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out9_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out10_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out10_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out11_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out11_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out12_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out12_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out13_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out13_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out14_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out14_im;
	wire	[WORD_SIZE-1:0]	w_buffer_out15_re;
	wire	[WORD_SIZE-1:0]	w_buffer_out15_im;	
	
	control_unit_FFT32	my_control_unit_FFT32
	(
		.i_clk(i_clk),
		.i_rst(i_rst),
		.w_FFT16_cycle_done(w_FFT16_cycle_done),
	
		.o_mux_switcher(w_mux_switcher),
		.o_address_switcher(w_address_switcher),
		.o_FFT16_cycle_rst(w_FFT16_cycle_rst),
		.o_STAGES(w_STAGES),
		.o_FFT16_cycle_done_delay(w_FFT16_cycle_done_delay),
		.o_FFT32_cycle_done(o_FFT32_cycle_done)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in0 
	(
		.a_re(in0_re),
		.a_im(in0_im),
		.b_re(in1_re),
		.b_im(in1_im),
		.c_re(out0_re),
		.c_im(out0_im),
		.d_re(w_buffer_out1_re),
		.d_im(w_buffer_out1_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in0_re),
		.out_im(FFT16_in0_im)
	);

	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in1 
	(
		.a_re(in2_re),
		.a_im(in2_im),
		.b_re(in3_re),
		.b_im(in3_im),
		.c_re(out8_re),
		.c_im(out8_im),
		.d_re(w_buffer_out9_re),
		.d_im(w_buffer_out9_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in1_re),
		.out_im(FFT16_in1_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in2 
	(
		.a_re(in4_re),
		.a_im(in4_im),
		.b_re(in5_re),
		.b_im(in5_im),
		.c_re(out4_re),
		.c_im(out4_im),
		.d_re(w_buffer_out5_re),
		.d_im(w_buffer_out5_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in2_re),
		.out_im(FFT16_in2_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in3 
	(
		.a_re(in6_re),
		.a_im(in6_im),
		.b_re(in7_re),
		.b_im(in7_im),
		.c_re(out12_re),
		.c_im(out12_im),
		.d_re(w_buffer_out13_re),
		.d_im(w_buffer_out13_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in3_re),
		.out_im(FFT16_in3_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in4 
	(
		.a_re(in8_re),
		.a_im(in8_im),
		.b_re(in9_re),
		.b_im(in9_im),
		.c_re(out2_re), 
		.c_im(out2_im), 
		.d_re(w_buffer_out3_re),
		.d_im(w_buffer_out3_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in4_re),
		.out_im(FFT16_in4_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in5 
	(
		.a_re(in10_re),
		.a_im(in10_im),
		.b_re(in11_re),
		.b_im(in11_im),
		.c_re(out10_re),
		.c_im(out10_im),
		.d_re(w_buffer_out11_re),
		.d_im(w_buffer_out11_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in5_re),
		.out_im(FFT16_in5_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in6 
	(
		.a_re(in12_re),
		.a_im(in12_im),
		.b_re(in13_re),
		.b_im(in13_im),
		.c_re(out6_re),
		.c_im(out6_im),
		.d_re(w_buffer_out7_re),
		.d_im(w_buffer_out7_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in6_re),
		.out_im(FFT16_in6_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in7 
	(
		.a_re(in14_re),
		.a_im(in14_im),
		.b_re(in15_re),
		.b_im(in15_im),
		.c_re(out14_re),
		.c_im(out14_im),
		.d_re(w_buffer_out15_re),
		.d_im(w_buffer_out15_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in7_re),
		.out_im(FFT16_in7_im)
	);
	
		mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in8 
	(
		.a_re(in16_re),
		.a_im(in16_im),
		.b_re(in17_re),
		.b_im(in17_im),
		.c_re(out16_re),
		.c_im(out16_im),
		.d_re(out17_re),
		.d_im(out17_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in8_re),
		.out_im(FFT16_in8_im)
	);

	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in9 
	(
		.a_re(in18_re),
		.a_im(in18_im),
		.b_re(in19_re),
		.b_im(in19_im),
		.c_re(out24_re),
		.c_im(out24_im),
		.d_re(out25_re),
		.d_im(out25_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in9_re),
		.out_im(FFT16_in9_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in10 
	(
		.a_re(in20_re),
		.a_im(in20_im),
		.b_re(in21_re),
		.b_im(in21_im),
		.c_re(out20_re),
		.c_im(out20_im),
		.d_re(out21_re),
		.d_im(out21_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in10_re),
		.out_im(FFT16_in10_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in11 
	(
		.a_re(in22_re),
		.a_im(in22_im),
		.b_re(in23_re),
		.b_im(in23_im),
		.c_re(out28_re),
		.c_im(out28_im),
		.d_re(out29_re),
		.d_im(out29_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in11_re),
		.out_im(FFT16_in11_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in12 
	(
		.a_re(in24_re),
		.a_im(in24_im),
		.b_re(in25_re),
		.b_im(in25_im),
		.c_re(out18_re), 
		.c_im(out18_im), 
		.d_re(out19_re),
		.d_im(out19_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in12_re),
		.out_im(FFT16_in12_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in13 
	(
		.a_re(in26_re),
		.a_im(in26_im),
		.b_re(in27_re),
		.b_im(in27_im),
		.c_re(out26_re),
		.c_im(out26_im),
		.d_re(out27_re),
		.d_im(out27_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in13_re),
		.out_im(FFT16_in13_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in14 
	(
		.a_re(in28_re),
		.a_im(in28_im),
		.b_re(in29_re),
		.b_im(in29_im),
		.c_re(out22_re),
		.c_im(out22_im),
		.d_re(out23_re),
		.d_im(out23_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in14_re),
		.out_im(FFT16_in14_im)
	);
	
	mux4in1_complex #(.WORD_SIZE(WORD_SIZE)) mux_FFT16_in15 
	(
		.a_re(in30_re),
		.a_im(in30_im),
		.b_re(in31_re),
		.b_im(in31_im),
		.c_re(out30_re),
		.c_im(out30_im),
		.d_re(out31_re),
		.d_im(out31_im),
		.sel(w_mux_switcher),
		.out_re(FFT16_in15_re),
		.out_im(FFT16_in15_im)
	);
	
	FFT16_top #(.WORD_SIZE(WORD_SIZE), .FRACTION(FRACTION)) FFT16
	(
		.i_clk(i_clk),
		.i_rst(w_FFT16_cycle_rst | i_rst),
		.STAGES(w_STAGES),
		.choose_twiddle(w_mux_switcher),
		.in0_re(FFT16_in0_re),
		.in0_im(FFT16_in0_im),
		.in1_re(FFT16_in1_re),
		.in1_im(FFT16_in1_im),
		.in2_re(FFT16_in2_re),
		.in2_im(FFT16_in2_im),
		.in3_re(FFT16_in3_re),
		.in3_im(FFT16_in3_im),
		.in4_re(FFT16_in4_re),
		.in4_im(FFT16_in4_im),
		.in5_re(FFT16_in5_re),
		.in5_im(FFT16_in5_im),
		.in6_re(FFT16_in6_re),
		.in6_im(FFT16_in6_im),
		.in7_re(FFT16_in7_re),
		.in7_im(FFT16_in7_im),
		.in8_re(FFT16_in8_re),
		.in8_im(FFT16_in8_im),
		.in9_re(FFT16_in9_re),
		.in9_im(FFT16_in9_im),
		.in10_re(FFT16_in10_re),
		.in10_im(FFT16_in10_im),
		.in11_re(FFT16_in11_re),
		.in11_im(FFT16_in11_im),
		.in12_re(FFT16_in12_re),
		.in12_im(FFT16_in12_im),
		.in13_re(FFT16_in13_re),
		.in13_im(FFT16_in13_im),
		.in14_re(FFT16_in14_re),
		.in14_im(FFT16_in14_im),
		.in15_re(FFT16_in15_re),
		.in15_im(FFT16_in15_im),
		
		.out0_re(FFT16_out0_re),
		.out0_im(FFT16_out0_im),
		.out1_re(FFT16_out1_re),
		.out1_im(FFT16_out1_im),
		.out2_re(FFT16_out2_re),
		.out2_im(FFT16_out2_im),
		.out3_re(FFT16_out3_re),
		.out3_im(FFT16_out3_im),
		.out4_re(FFT16_out4_re),
		.out4_im(FFT16_out4_im),
		.out5_re(FFT16_out5_re),
		.out5_im(FFT16_out5_im),
		.out6_re(FFT16_out6_re),
		.out6_im(FFT16_out6_im),
		.out7_re(FFT16_out7_re),
		.out7_im(FFT16_out7_im),
		.out8_re(FFT16_out8_re),
		.out8_im(FFT16_out8_im),
		.out9_re(FFT16_out9_re),
		.out9_im(FFT16_out9_im),
		.out10_re(FFT16_out10_re),
		.out10_im(FFT16_out10_im),
		.out11_re(FFT16_out11_re),
		.out11_im(FFT16_out11_im),
		.out12_re(FFT16_out12_re),
		.out12_im(FFT16_out12_im),
		.out13_re(FFT16_out13_re),
		.out13_im(FFT16_out13_im),
		.out14_re(FFT16_out14_re),
		.out14_im(FFT16_out14_im),
		.out15_re(FFT16_out15_re),
		.out15_im(FFT16_out15_im),

		.o_FFT_cycle_done(w_FFT16_cycle_done)
	);

	ram_16_byte #( .WORD_SIZE(WORD_SIZE)) buffer_ram
	(
		.we(w_FFT16_cycle_done_delay && ~w_address_switcher && (w_mux_switcher < 2)),
		.in0_re(FFT16_out0_re),
		.in0_im(FFT16_out0_im),
		.in1_re(FFT16_out1_re),
		.in1_im(FFT16_out1_im),
		.in2_re(FFT16_out2_re),
		.in2_im(FFT16_out2_im),
		.in3_re(FFT16_out3_re),
		.in3_im(FFT16_out3_im),
		.in4_re(FFT16_out4_re),
		.in4_im(FFT16_out4_im),
		.in5_re(FFT16_out5_re),
		.in5_im(FFT16_out5_im),
		.in6_re(FFT16_out6_re),
		.in6_im(FFT16_out6_im),
		.in7_re(FFT16_out7_re),
		.in7_im(FFT16_out7_im),
		.in8_re(FFT16_out8_re),
		.in8_im(FFT16_out8_im),
		.in9_re(FFT16_out9_re),
		.in9_im(FFT16_out9_im),
		.in10_re(FFT16_out10_re),
		.in10_im(FFT16_out10_im),
		.in11_re(FFT16_out11_re),
		.in11_im(FFT16_out11_im),
		.in12_re(FFT16_out12_re),
		.in12_im(FFT16_out12_im),
		.in13_re(FFT16_out13_re),
		.in13_im(FFT16_out13_im),
		.in14_re(FFT16_out14_re),
		.in14_im(FFT16_out14_im),
		.in15_re(FFT16_out15_re),
		.in15_im(FFT16_out15_im),
		
		.out0_re(w_buffer_out0_re),
		.out0_im(w_buffer_out0_im),
		.out1_re(w_buffer_out1_re),
		.out1_im(w_buffer_out1_im),
		.out2_re(w_buffer_out2_re),
		.out2_im(w_buffer_out2_im),
		.out3_re(w_buffer_out3_re),
		.out3_im(w_buffer_out3_im),
		.out4_re(w_buffer_out4_re),
		.out4_im(w_buffer_out4_im),
		.out5_re(w_buffer_out5_re),
		.out5_im(w_buffer_out5_im),
		.out6_re(w_buffer_out6_re),
		.out6_im(w_buffer_out6_im),
		.out7_re(w_buffer_out7_re),
		.out7_im(w_buffer_out7_im),
		.out8_re(w_buffer_out8_re),
		.out8_im(w_buffer_out8_im),
		.out9_re(w_buffer_out9_re),
		.out9_im(w_buffer_out9_im),
		.out10_re(w_buffer_out10_re),
		.out10_im(w_buffer_out10_im),
		.out11_re(w_buffer_out11_re),
		.out11_im(w_buffer_out11_im),
		.out12_re(w_buffer_out12_re),
		.out12_im(w_buffer_out12_im),
		.out13_re(w_buffer_out13_re),
		.out13_im(w_buffer_out13_im),
		.out14_re(w_buffer_out14_re),
		.out14_im(w_buffer_out14_im),
		.out15_re(w_buffer_out15_re),
		.out15_im(w_buffer_out15_im)
	);

	ram_32_byte #(.WORD_SIZE(WORD_SIZE)) my_ram_32_byte 
	(
		.we(w_FFT16_cycle_done_delay),
		.address(w_address_switcher),
		.in0_re(FFT16_out0_re),
		.in0_im(FFT16_out0_im),
		.in1_re(FFT16_out1_re),
		.in1_im(FFT16_out1_im),
		.in2_re(FFT16_out2_re),
		.in2_im(FFT16_out2_im),
		.in3_re(FFT16_out3_re),
		.in3_im(FFT16_out3_im),
		.in4_re(FFT16_out4_re),
		.in4_im(FFT16_out4_im),
		.in5_re(FFT16_out5_re),
		.in5_im(FFT16_out5_im),
		.in6_re(FFT16_out6_re),
		.in6_im(FFT16_out6_im),
		.in7_re(FFT16_out7_re),
		.in7_im(FFT16_out7_im),
		.in8_re(FFT16_out8_re),
		.in8_im(FFT16_out8_im),
		.in9_re(FFT16_out9_re),
		.in9_im(FFT16_out9_im),
		.in10_re(FFT16_out10_re),
		.in10_im(FFT16_out10_im),
		.in11_re(FFT16_out11_re),
		.in11_im(FFT16_out11_im),
		.in12_re(FFT16_out12_re),
		.in12_im(FFT16_out12_im),
		.in13_re(FFT16_out13_re),
		.in13_im(FFT16_out13_im),
		.in14_re(FFT16_out14_re),
		.in14_im(FFT16_out14_im),
		.in15_re(FFT16_out15_re),
		.in15_im(FFT16_out15_im),
		
		.out0_re(out0_re),
		.out0_im(out0_im),
		.out1_re(out1_re),
		.out1_im(out1_im),
		.out2_re(out2_re),
		.out2_im(out2_im),
		.out3_re(out3_re),
		.out3_im(out3_im),
		.out4_re(out4_re),
		.out4_im(out4_im),
		.out5_re(out5_re),
		.out5_im(out5_im),
		.out6_re(out6_re),
		.out6_im(out6_im),
		.out7_re(out7_re),
		.out7_im(out7_im),
		.out8_re(out8_re),
		.out8_im(out8_im),
		.out9_re(out9_re),
		.out9_im(out9_im),
		.out10_re(out10_re),
		.out10_im(out10_im),
		.out11_re(out11_re),
		.out11_im(out11_im),
		.out12_re(out12_re),
		.out12_im(out12_im),
		.out13_re(out13_re),
		.out13_im(out13_im),
		.out14_re(out14_re),
		.out14_im(out14_im),
		.out15_re(out15_re),
		.out15_im(out15_im),
		.out16_re(out16_re),
		.out16_im(out16_im),
		.out17_re(out17_re),
		.out17_im(out17_im),
		.out18_re(out18_re),
		.out18_im(out18_im),
		.out19_re(out19_re),
		.out19_im(out19_im),
		.out20_re(out20_re),
		.out20_im(out20_im),
		.out21_re(out21_re),
		.out21_im(out21_im),
		.out22_re(out22_re),
		.out22_im(out22_im),
		.out23_re(out23_re),
		.out23_im(out23_im),
		.out24_re(out24_re),
		.out24_im(out24_im),
		.out25_re(out25_re),
		.out25_im(out25_im),
		.out26_re(out26_re),
		.out26_im(out26_im),
		.out27_re(out27_re),
		.out27_im(out27_im),
		.out28_re(out28_re),
		.out28_im(out28_im),
		.out29_re(out29_re),
		.out29_im(out29_im),
		.out30_re(out30_re),
		.out30_im(out30_im),
		.out31_re(out31_re),
		.out31_im(out31_im)
	);

endmodule