module mux32in1 #(parameter DATA_LENGTH = 8)
(
	input 	[DATA_LENGTH-1:0]		in1,
	input 	[DATA_LENGTH-1:0]		in2,
	input 	[DATA_LENGTH-1:0]		in3,
	input 	[DATA_LENGTH-1:0]		in4,
	input 	[DATA_LENGTH-1:0]		in5,
	input 	[DATA_LENGTH-1:0]		in6,
	input 	[DATA_LENGTH-1:0]		in7,
	input 	[DATA_LENGTH-1:0]		in8,
	input 	[DATA_LENGTH-1:0]		in9,
	input 	[DATA_LENGTH-1:0]		in10
);


endmodule
